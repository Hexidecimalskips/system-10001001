��1   1 0   1 1   1 0 0   1 0 1   1 1 0   1 1 1   1 0 0 0   1 0 0 1   1 0 1 0   1 0 1 1   1 1 0 0   1 1 0 1   1 1 1 0   1 1 1 1   1 0 0 0 0   1 0 0 0 1   1 0 0 1 0   1 0 0 1 1   1 0 1 0 0   1 0 1 0 1   1 0 1 1 0   1 0 1 1 1   1 1 0 0 0   1 1 0 0 1   1 1 0 1 0   1 1 0 1 1   1 1 1 0 0   1 1 1 0 1   1 1 1 1 0   1 1 1 1 1   1 0 0 0 0 0   1 0 0 0 0 1   1 0 0 0 1 0   1 0 0 0 1 1   1 0 0 1 0 1   1 0 0 1 1 0   1 0 0 1 1 1   1 0 1 0 0 0   1 0 1 0 0 1   1 0 1 0 1 0   1 0 1 0 1 1   1 0 1 1 0 0   1 0 1 1 0 1   1 0 1 1 1 0   1 0 1 1 1 1   1 1 0 0 0 0   1 1 0 0 0 1   1 1 0 0 1 0   1 1 0 0 1 1   1 1 0 1 0 0   1 1 0 1 0 1   1 1 0 1 1 0   1 1 0 1 1 1   1 1 1 0 0 0   1 1 1 0 0 1   1 1 1 0 1 0   1 1 1 0 1 1   1 1 1 1 0 0   1 1 1 1 0 1   1 1 1 1 1 0   1 1 1 1 1 1   1 0 0 0 0 0 0   1 0 0 0 0 0 1   1 0 0 0 0 1 0   1 0 0 0 0 1 1   1 0 0 0 1 0 0   1 0 0 0 1 0 1   1 0 0 0 1 1 0   1 0 0 0 1 1 1   1 0 0 1 0 0 0   1 0 0 1 0 0 1   1 0 0 1 0 1 0   1 0 0 1 0 1 1   1 0 0 1 1 0 0   1 0 0 1 1 0 1   1 0 0 1 1 1 0   1 0 0 1 1 1 1   1 0 1 0 0 0 0   1 0 1 0 0 0 1   1 0 1 0 0 1 0   1 0 1 0 0 1 1   1 0 1 0 1 0 0   1 0 1 0 1 0 1   1 0 1 0 1 1 0   1 0 1 0 1 1 1   1 0 1 1 0 0 0   1 0 1 1 0 0 1   1 0 1 1 0 1 0   1 0 1 1 0 1 1   1 0 1 1 1 0 0   1 0 1 1 1 0 1   1 0 1 1 1 1 0   1 0 1 1 1 1 1   1 1 0 0 0 0 0   1 1 1 0 0 0 0   1 1 1 0 0 0 1   1 1 1 1 0 0 0   1 1 1 1 0 0 1   1 1 1 1 0 1 0   1 1 1 1 0 1 1   1 1 1 1 1 0 0   1 1 1 1 1 0 1   1 1 1 1 1 1 0   1 1 1 1 1 1 1   1 0 0 0 0 0 0 0   1 0 0 0 0 0 0 1   1 0 0 0 0 0 1 0   1 0 0 0 0 0 1 1   1 0 0 0 0 1 0 0   1 0 0 0 0 1 0 1   1 0 0 0 0 1 1 0   1 0 0 0 0 1 1 1   1 0 0 0 1 0 0 0   1 0 0 1 0 0 0 1   1 0 0 0 1 0 1 1   1 0 0 0 1 1 0 1   1 0 0 0 1 1 1 0   1 0 0 0 1 1 1 1   1 0 0 1 0 0 0 0   1 0 0 1 0 0 0 1   1 0 0 1 0 0 1 0   1 0 0 1 0 0 1 1   1 0 0 1 0 1 0 0   1 0 0 1 0 1 0 1   1 0 0 1 0 1 1 0   1 0 0 1 0 1 1 1   1 0 0 1 1 0 0 0   1 0 0 1 1 0 0 1   1 0 0 1 1 0 1 0   1 0 0 1 1 0 1 1   1 0 0 1 1 1 0 0   1 0 0 1 1 1 0 1   1 0 0 1 1 1 1 0   1 0 0 1 1 1 1 1   1 0 1 0 0 0 0 0   1 0 1 0 0 0 0 1   1 0 1 0 0 0 1 0   1 0 1 0 0 0 1 1   1 0 1 0 0 1 0 0   1 0 1 0 0 1 0 1   1 0 1 0 0 1 1 0   1 0 1 0 0 1 1 1   1 0 1 0 1 0 0 0   1 0 1 0 1 0 0 1   1 0 1 0 1 0 1 0   1 0 1 0 1 0 1 1   1 0 1 0 1 1 0 0   1 0 1 0 1 1 0 1   1 0 1 0 1 1 1 0   1 0 1 0 1 1 1 1   1 0 1 1 0 0 0 0   1 0 1 1 0 0 0 1   1 0 1 1 0 0 1 0   1 0 1 1 0 0 1 1   1 0 1 1 0 1 0 0   1 0 1 1 0 1 0 1   1 0 1 1 0 1 1 0   1 0 1 1 0 1 1 1   1 0 1 1 1 0 0 0   1 0 1 1 1 0 0 1   1 0 1 1 1 0 1 0   1 0 1 1 1 0 1 1   1 0 1 1 1 1 0 0   1 0 1 1 1 1 0 1   1 0 1 1 1 1 1 0   1 0 1 1 1 1 1 1   1 1 0 0 0 0 0 0   1 1 0 0 0 0 0 1   1 1 0 0 0 0 1 0   1 1 0 0 0 0 1 1   1 1 0 0 0 1 0 0   1 1 0 0 0 1 0 1   1 1 0 0 0 1 1 0   1 1 0 0 0 1 1 1   1 1 0 0 1 0 0 0   1 1 0 0 1 0 0 1   1 1 0 0 1 0 1 0   1 1 0 0 1 0 1 1   1 1 0 0 1 1 0 0   1 1 0 0 1 1 0 1   1 1 0 0 1 1 1 0   1 1 0 0 1 1 1 1   1 1 0 1 0 0 0 0   1 1 0 1 0 0 0 1   1 1 0 1 0 0 1 0   1 1 0 1 0 0 1 1   1 1 0 1 0 1 0 0   1 1 0 1 0 1 0 1   1 1 0 1 0 1 1 0   1 1 0 1 0 1 1 1   1 1 0 1 1 0 0 0   1 1 0 1 1 0 0 1   1 1 0 1 1 0 1 0   1 1 0 1 1 0 1 1   1 1 0 1 1 1 0 0   1 1 0 1 1 1 0 1   1 1 0 1 1 1 1 0   1 1 0 1 1 1 1 1   1 1 1 0 0 0 0 0   1 1 1 0 0 0 0 1   1 1 1 0 0 0 1 0   1 1 1 0 0 0 1 1   1 1 1 0 0 1 0 0   1 1 1 0 0 1 0 1   1 1 1 0 0 1 1 0   1 1 1 0 0 1 1 1   1 1 1 0 1 0 0 0   1 1 1 0 1 0 0 1   1 1 1 0 1 0 1 0   1 1 1 0 1 0 1 1   1 1 1 0 1 1 0 0   1 1 1 0 1 1 0 1   1 1 1 0 1 1 1 0   1 1 1 0 1 1 1 1   1 1 1 1 0 0 0 0   1 1 1 1 0 0 0 1   1 1 1 1 0 0 1 0   1 1 1 1 0 0 1 1   1 1 1 1 0 1 0 0   1 1 1 1 0 1 0 1   1 1 1 1 0 1 1 0   1 1 1 1 1 0 0 0   1 1 1 1 1 0 0 1   1 1 1 1 1 0 1 0   1 1 1 1 1 0 1 1   1 1 1 1 1 1 0 0   1 1 1 1 1 1 0 1   1 1 1 1 1 1 1 0   1 1 1 1 1 1 1 1   1 1 1 1 1 1 1 0   1 1 1 1 1 1 0 1   1 1 1 1 1 1 0 0   1 1 1 1 1 0 1 1   1 1 1 1 1 0 1 0   1 1 1 1 1 0 0 1   1 1 1 1 1 0 0 0   1 1 1 1 0 1 1 1   1 1 1 1 0 1 1 0   1 1 1 1 0 1 0 1   1 1 1 1 0 1 0 0   1 1 1 1 0 0 1 1   1 1 1 1 0 0 1 0   1 1 1 1 0 0 0 1   1 1 1 1 0 0 0 0   1 1 1 0 1 1 1 1   1 1 1 0 1 1 1 0   1 1 1 0 1 1 0 1   1 1 1 0 1 1 0 0   1 1 1 0 1 0 1 1   1 1 1 0 1 0 1 0   1 1 1 0 1 0 0 1   1 1 1 0 1 0 0 0   1 1 1 0 0 1 1 1   1 1 1 0 0 1 1 0   1 1 1 0 0 1 0 1   1 1 1 0 0 1 0 0   1 1 1 0 0 0 1 1   1 1 1 0 0 0 1 0   1 1 1 0 0 0 0 1   1 1 1 0 0 0 0 0   1 1 0 1 1 1 1 0   1 1 0 1 1 1 0 1   1 1 0 1 1 1 0 0   1 1 0 1 1 0 1 1   1 1 0 1 1 0 1 0   1 1 0 1 1 0 0 1   1 1 0 1 1 0 0 0   1 1 0 1 0 1 1 1   1 1 0 1 0 1 1 0   1 1 0 1 0 1 0 1   1 1 0 1 0 1 0 0   1 1 0 1 0 0 1 1   1 1 0 1 0 0 1 0   1 1 0 1 0 0 0 1   1 1 0 1 0 0 0 0   1 1 0 0 1 1 1 1   1 1 0 0 1 1 1 0   1 1 0 0 1 1 0 1   1 1 0 0 1 1 0 0   1 1 0 0 1 0 1 1   1 1 0 0 1 0 1 0   1 1 0 0 1 0 0 1   1 1 0 0 1 0 0 0   1 1 0 0 0 1 1 1   1 1 0 0 0 1 1 0   1 1 0 0 0 1 0 1   1 1 0 0 0 1 0 0   1 1 0 0 0 0 1 1   1 1 0 0 0 0 1 0   1 1 0 0 0 0 0 1   1 1 0 0 0 0 0 0   1 0 1 1 1 1 1 0   1 0 1 1 1 1 0 1   1 0 1 1 1 1 0 0   1 0 1 1 1 0 1 1   1 0 1 1 1 0 1 0   1 0 1 1 1 0 0 1   1 0 1 1 1 0 0 0   1 0 1 1 0 1 1 1   1 0 1 1 0 1 1 0   1 0 1 1 0 1 0 1   1 0 1 1 0 1 0 0   1 0 1 1 0 0 1 1   1 0 1 1 0 0 1 0   1 0 1 1 0 0 0 1   1 0 1 1 0 0 0 0   1 0 1 0 1 1 1 1   1 0 1 0 1 1 1 0   1 0 1 0 1 1 0 1   1 0 1 0 1 1 0 0   1 0 1 0 1 0 1 1   1 0 1 0 1 0 1 0   1 0 1 0 1 0 0 1   1 0 1 0 1 0 0 0   1 0 1 0 0 1 1 1   1 0 1 0 0 1 1 0   1 0 1 0 0 1 0 1   1 0 1 0 0 1 0 0   1 0 1 0 0 0 1 1   1 0 1 0 0 0 1 0   1 0 1 0 0 0 0 1   1 0 1 0 0 0 0 0   1 0 0 1 1 1 1 0   1 0 0 1 1 1 0 1   1 0 0 1 1 1 0 0   1 0 0 1 1 0 1 1   1 0 0 1 1 0 1 0   1 0 0 1 1 0 0 1   1 0 0 1 1 0 0 0   1 0 0 1 0 1 1 1   1 0 0 1 0 1 1 0   1 0 0 1 0 1 0 1   1 0 0 1 0 1 0 0   1 0 0 1 0 0 1 1   1 0 0 1 0 0 1 0   1 0 0 1 0 0 0 1   1 0 0 1 0 0 0 0   1 0 0 0 1 1 1 1   1 0 0 0 1 1 1 0   1 0 0 0 1 1 0 1   1 0 0 0 1 1 0 0   1 0 0 0 1 0 1 1   1 0 0 0 1 0 1 0   1 0 0 0 1 0 0 1   1 0 0 0 1 0 0 0   1 0 0 0 0 1 1 1   1 0 0 0 0 1 1 0   1 0 0 0 0 1 0 1   1 0 0 0 0 1 0 0   1 0 0 0 0 0 1 1   1 0 0 0 0 0 1 0   1 0 0 0 0 0 0 1   1 0 0 0 0 0 0 0   0 1 1 1 1 1 1 0   0 1 1 1 1 1 0 1   0 1 1 1 1 1 0 0   0 1 1 1 1 0 1 1   0 1 1 1 1 0 1 0   0 1 1 1 1 0 0 1   0 1 1 1 1 0 0 0   0 1 1 1 0 1 1 1   0 1 1 1 0 1 1 0   0 1 1 1 0 1 0 1   0 1 1 1 0 1 0 0   0 1 1 1 0 0 1 1   0 1 1 1 0 0 1 0   0 1 1 1 0 0 0 1   0 1 1 1 0 0 0 0   0 1 1 0 1 1 1 1   0 1 1 0 1 1 1 0   0 1 1 0 1 1 0 1   0 1 1 0 1 1 0 0   0 1 1 0 1 0 1 1   0 1 1 0 1 0 1 0   0 1 1 0 1 0 0 1   0 1 1 0 1 0 0 0   0 1 1 0 0 1 1 1   0 1 1 0 0 1 1 0   0 1 1 0 0 1 0 1   0 1 1 0 0 1 0 0   0 1 1 0 0 0 1 1   0 1 1 0 0 0 0 1   0 1 1 0 0 0 0 0   0 1 0 1 1 1 1 1   0 1 0 1 1 1 1 0   0 1 0 1 1 1 0 1   0 1 0 1 1 1 0 0   0 1 0 1 1 0 1 1   0 1 0 1 1 0 1 0   0 1 0 1 1 0 0 1   0 1 0 1 1 0 0 0   0 1 0 1 0 1 1 1   0 1 0 1 0 1 1 0   0 1 0 1 0 1 0 1   0 1 0 1 0 1 0 0   0 1 0 1 0 0 1 1   0 1 0 1 0 0 1 0   0 1 0 1 0 0 0 1   0 1 0 1 0 0 0 0   0 1 0 0 1 1 1 0   0 1 0 0 1 1 0 1   0 1 0 0 1 1 0 0   0 1 0 0 1 0 1 1   0 1 0 0 1 0 1 0   0 1 0 0 1 0 0 1   0 1 0 0 1 0 0 0   0 1 0 0 0 1 1 1   0 1 0 0 0 1 1 0   0 1 0 0 0 1 0 1   0 1 0 0 0 1 0 0   0 1 0 0 0 0 1 1   0 1 0 0 0 0 1 0   0 1 0 0 0 0 0 1   0 1 0 0 0 0 0 0   0 0 1 1 1 1 1 0   0 0 1 1 1 1 0 1   0 0 1 1 1 1 0 0   0 0 1 1 1 0 1 1   0 0 1 1 1 0 1 0   0 0 1 1 1 0 0 1   0 0 1 1 1 0 0 0   0 0 1 1 0 1 1 1   0 0 1 1 0 1 1 0   0 0 1 1 0 1 0 1   0 0 1 1 0 1 0 0   0 0 1 1 0 0 1 1   0 0 1 1 0 0 1 0   0 0 1 1 0 0 0 1   0 0 1 1 0 0 0 0   0 0 1 0 1 1 1 1   0 0 1 0 1 1 1 0   0 0 1 0 1 1 0 1   0 0 1 0 1 1 0 0   0 0 1 0 1 0 1 1   0 0 1 0 1 0 1 0   0 0 1 1 0 0 0 1   0 0 1 0 1 0 1 0   0 0 1 0 1 0 0 1   0 0 1 0 1 0 0 0   0 0 1 0 0 1 1 1   0 0 1 0 0 1 1 0   0 0 1 0 0 1 0 1   0 0 1 0 0 1 0 0   0 0 1 0 0 0 1 1   0 0 1 0 0 0 1 0   0 0 1 0 0 0 0 1   0 0 1 0 0 0 0 0   0 0 0 1 1 1 1 1   0 0 0 0 1 1 1 1   0 0 0 0 1 1 1 0   0 0 0 0 1 1 0 1   0 0 0 0 1 1 0 0   0 0 0 0 1 0 1 1   0 0 0 0 1 0 1 0   0 0 0 0 1 0 0 1   0 0 0 0 1 0 0 0   0 0 0 0 0 1 1 1   0 0 0 0 0 1 1 0   0 0 0 0 0 1 0 1   0 0 0 0 0 1 0 0   0 0 0 0 0 0 1 1   0 0 0 0 0 0 1 0   0 0 0 0 0 0 0 1   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0   0 0 0 0 0 0 0     0 0 0 0 0 0 0 0     0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   3 : 2 3   P M   2 0 2 4 - 1 2 - 2 6  
 1 0 0 0 0 0 0 0 1   1 0 0 0 1 0 0 0 1   1 0 0 0 1 0 0 1 0   1 0 0 0 1 0 0 1 1   1 0 0 0 1 0 1 0 0   1 0 0 0 1 0 1 0 1   1 0 0 0 1 0 1 1 0   1 0 0 0 1 0 1 1 1   1 0 0 0 1 1 0 0 0   1 0 0 0 1 1 0 0 1   1 0 0 0 1 1 0 1 0   1 0 0 0 1 1 0 1 1   1 0 0 0 1 1 1 0 0   1 0 0 0 1 1 1 0 1   1 0 0 0 1 1 1 1 0   1 0 0 0 1 1 1 1 1   1 0 0 1 0 0 0 0 0   1 0 0 1 0 0 0 0 1   1 0 0 1 0 0 0 1 0   1 0 0 1 0 0 0 1 1   1 0 0 1 0 0 1 0 0   1 0 0 1 0 0 1 0 1   1 0 0 1 0 0 1 1 0   1 0 0 1 0 0 1 1 1   1 0 0 1 0 1 0 0 0   1 0 0 1 0 1 0 0 1   1 0 0 1 0 1 0 1 0   1 0 0 1 0 1 0 1 1   1 0 0 1 0 1 1 0 0   1 0 0 1 0 1 1 0 1   1 0 0 1 0 1 1 1 0   1 0 0 1 0 1 1 1 1   1 0 0 1 1 0 0 0 0   1 0 0 1 1 0 0 0 1   1 0 0 1 1 0 0 1 0   1 0 0 1 1 0 0 1 1   1 0 0 1 1 0 1 0 0   1 0 0 1 1 0 1 0 1   1 0 0 1 1 0 1 1 0   1 0 0 1 1 0 1 1 1   1 0 0 1 1 1 0 0 0   1 0 0 1 1 1 0 0 1   1 0 0 1 1 1 0 0 1   1 0 0 1 1 1 0 1 0   1 0 0 1 1 1 0 1 1   1 0 0 1 1 1 1 0 0   1 0 0 1 1 1 1 0 1   1 0 0 1 1 1 1 1 0   1 0 0 1 1 1 1 1 1   1 0 1 0 0 0 0 0 0   1 0 1 0 0 0 0 0 1   1 0 1 0 0 0 0 1 0   1 0 1 0 0 0 0 1 1   1 0 1 0 0 0 1 0 0   1 0 1 0 0 0 1 0 1   1 0 1 0 0 0 1 1 0   1 0 1 0 0 0 1 1 1   1 0 1 0 0 1 0 0 0   1 0 1 0 0 1 0 0 1   1 0 1 0 0 1 0 1 0   1 0 1 0 0 1 0 1 1   1 0 1 0 0 1 1 0 0   1 0 1 0 0 1 1 0 1   1 0 1 0 0 1 1 1 0   1 0 1 0 0 1 1 1 1   1 0 1 0 1 0 0 0 0   1 0 1 0 1 0 0 0 1   1 0 1 0 1 0 0 1 0   1 0 1 0 1 0 0 1 1   1 0 1 0 1 0 1 0 0   1 0 1 0 1 0 1 0 1   1 0 1 0 1 0 1 1 0   1 0 1 0 1 0 1 1 1   1 0 1 0 1 1 0 0 0   1 0 1 0 1 1 0 0 1   1 0 1 0 1 1 0 1 0   1 0 1 0 1 1 0 1 1   1 0 1 0 1 1 1 0 0   1 0 1 0 1 1 1 0 1   1 0 1 0 1 1 1 1 0   1 0 1 0 1 1 1 1 1   1 0 1 1 0 0 0 0 0   1 0 1 1 0 0 0 0 1   1 0 1 1 0 0 0 1 0   1 0 1 1 0 0 0 1 1   1 0 1 1 0 0 1 0 0   1 0 1 1 0 0 1 0 1   1 0 1 1 0 0 1 1 0   1 0 1 1 0 0 1 1 1   1 0 1 1 0 1 0 0 0   1 0 1 1 0 1 0 0 1   1 0 1 1 0 1 0 1 0   1 0 1 1 0 1 0 1 1   1 0 1 1 0 1 1 0 0   1 0 1 1 0 1 1 0 1   1 0 1 1 0 1 1 1 0   1 0 1 1 0 1 1 1 1   1 0 1 1 1 0 0 0 0   1 0 1 1 1 0 0 0 1   1 0 1 1 1 0 0 1 0   1 0 1 1 1 0 0 1 1   1 0 1 1 1 0 1 0 0   1 0 1 1 1 0 1 0 1   1 0 1 1 1 0 1 1 0   1 0 1 1 1 0 1 1 1   1 0 1 1 1 1 0 0 0   1 0 1 1 1 1 0 0 1   1 0 1 1 1 1 0 1 0   1 0 1 1 1 1 0 1 1   1 0 1 1 1 1 1 0 0   1 0 1 1 1 1 1 0 1   1 0 1 1 1 1 1 1 0   1 0 1 1 1 1 1 1 1   1 1 0 0 0 0 0 0 0   1 1 0 0 0 0 0 0 1   1 1 0 0 0 0 0 1 0   1 1 0 0 0 0 0 1 1   1 1 0 0 0 0 1 0 0   1 1 0 0 0 0 1 0 1   1 1 0 0 0 0 1 1 0   1 1 0 0 0 0 1 1 1   1 1 0 0 0 1 0 0 0   1 1 0 0 0 1 0 0 1   1 1 0 0 0 1 0 1 0   1 1 0 0 0 1 0 1 1   1 1 0 0 0 1 1 0 0   1 1 0 0 0 1 1 0 1   1 1 0 0 0 1 1 1 0   1 1 0 0 0 1 1 1 1   1 1 0 0 1 0 0 0 0   1 1 0 0 1 0 0 0 1   1 1 0 0 1 0 0 1 0   1 1 0 0 1 0 0 1 1   1 1 0 0 1 0 1 0 0   1 1 0 0 1 0 1 0 1   1 1 0 0 1 0 1 1 0   1 1 0 0 1 0 1 1 1   1 1 0 0 1 1 0 0 0   1 1 0 0 1 1 0 0 1   1 1 0 0 1 1 0 1 0   1 1 0 0 1 1 0 1 1   1 1 0 0 1 1 1 0 0   1 1 0 0 1 1 1 0 1   1 1 0 0 1 1 1 1 0   1 1 0 0 1 1 1 1 1   1 1 0 1 0 0 0 0 0   1 1 0 1 0 0 0 0 1   1 1 0 1 0 0 0 1 0   1 1 0 1 0 0 0 1 1   1 1 0 1 0 0 1 0 0   1 1 0 1 0 0 1 0 1   1 1 0 1 0 0 1 1 0   1 1 0 1 0 0 1 1 1   1 1 0 1 0 1 0 0 0   1 1 0 1 0 1 0 0 1   1 1 0 1 0 1 0 1 0   1 1 0 1 0 1 0 1 1   1 1 0 1 0 1 1 0 0   1 1 0 1 0 1 1 0 1   1 1 0 1 0 1 1 1 0   1 1 0 1 0 1 1 1 1   1 1 0 1 1 0 0 0 0   1 1 0 1 1 0 0 0 1   1 1 0 1 1 0 0 1 0   1 1 0 1 1 0 0 1 1   1 1 0 1 1 0 1 0 0   1 1 0 1 1 0 1 0 1   1 1 0 1 1 0 1 1 0   1 1 0 1 1 0 1 1 1   1 1 0 1 1 1 0 0 0   1 1 0 1 1 1 0 0 1   1 1 0 1 1 1 0 1 0   1 1 0 1 1 1 0 1 1   1 1 0 1 1 1 1 0 0   1 1 0 1 1 1 0 1 1   1 1 0 1 1 1 1 0 1   1 1 0 1 1 1 1 1 0   1 1 0 1 1 1 1 1 1   1 1 1 0 0 0 0 0 0   1 1 1 0 0 0 0 0 1   1 1 1 0 0 0 0 1 0   1 1 1 0 0 0 0 1 1   1 1 1 0 0 0 1 0 0   1 1 1 0 0 0 1 0 1   1 1 1 0 0 0 1 1 0   1 1 1 0 0 0 1 1 1   1 1 1 0 0 1 0 0 0   1 1 1 0 0 1 0 0 1   1 1 1 0 0 1 0 1 0   1 1 1 0 0 1 0 1 1   1 1 1 0 0 1 1 0 0   1 1 1 0 0 1 1 0 1   1 1 1 0 0 1 1 1 0   1 1 1 0 0 1 1 1 1   1 1 1 0 1 0 0 0 0   1 1 1 0 1 0 0 0 1   1 1 1 0 1 0 0 1 0   1 1 1 0 1 0 0 1 1   1 1 1 0 1 0 1 0 0   1 1 1 0 1 0 1 0 1   1 1 1 0 1 0 1 1 0   1 1 1 0 1 0 1 1 1   1 1 1 0 1 1 0 0 0   1 1 1 0 1 1 0 0 1   1 1 1 0 1 1 0 1 0   1 1 1 0 1 1 0 1 1   1 1 1 0 1 1 1 0 0   1 1 1 0 1 1 1 0 1   1 1 1 0 1 1 1 1 0   1 1 1 0 1 1 1 1 1   1 1 1 1 0 0 0 0 0   1 1 1 1 0 0 0 0 1   1 1 1 1 0 0 0 1 0   1 1 1 1 0 0 0 1 1   1 1 1 1 0 0 1 0 0   1 1 1 1 0 0 1 0 1   1 1 1 1 0 0 1 1 0   1 1 1 1 0 0 1 1 1   1 1 1 1 0 1 0 0 0   1 1 1 1 0 1 0 0 1   1 1 1 1 0 1 0 1 0   1 1 1 1 0 1 0 1 1   1 1 1 1 0 1 1 0 0   1 1 1 1 0 1 1 0 1   1 1 1 1 0 1 1 1 0   1 1 1 1 0 1 1 1 1   1 1 1 1 1 0 0 0 0   1 1 1 1 1 0 0 0 1   1 1 1 1 1 0 0 1 0   1 1 1 1 1 0 0 1 1   1 1 1 1 1 0 1 0 0   1 1 1 1 1 0 1 0 1   1 1 1 1 1 0 1 1 0   1 1 1 1 1 0 1 1 1   1 1 1 1 1 1 0 0 0   1 1 1 1 1 1 0 0 1   1 1 1 1 1 1 0 1 0   1 1 1 1 1 1 0 1 1   1 1 1 1 1 1 0 0 0   1 1 1 1 1 1 0 0 1   1 1 1 1 1 1 0 1 0   1 1 1 1 1 1 0 1 1   1 1 1 1 1 1 1 0 0   1 1 1 1 1 1 1 0 1   1 1 1 1 1 1 1 1 0   1 1 1 1 1 1 1 1 1   1 1 1 1 1 1 1 1 0   1 1 1 1 1 1 1 0 1   1 1 1 1 1 1 1 0 0   1 1 1 1 1 1 0 1 1   1 1 1 1 1 1 0 1 0   1 1 1 1 1 1 0 0 1   1 1 1 1 1 1 0 0 0   1 1 1 1 1 0 1 1 1   1 1 1 1 1 0 1 1 0   1 1 1 1 1 0 1 0 1   1 1 1 1 1 0 1 0 0   1 1 1 1 1 0 0 1 1   1 1 1 1 1 0 0 0 1   1 1 1 1 1 0 0 0 0   1 1 1 1 0 1 1 1 1   1 1 1 1 0 1 1 1 0   1 1 1 1 0 1 1 0 1   1 1 1 1 0 1 1 0 0   1 1 1 1 0 1 0 1 1   1 1 1 1 0 1 0 1 0   1 1 1 1 0 1 0 0 1   1 1 1 1 0 1 0 0 0   1 1 1 1 0 0 1 1 1   1 1 1 1 0 0 1 1 0   1 1 1 1 0 0 1 0 1   1 1 1 1 0 0 1 0 0   1 1 1 1 0 0 0 1 1   1 1 1 1 0 0 0 1 0   1 1 1 1 0 0 0 0 1   1 1 1 1 0 0 0 0 0   1 1 1 0 1 1 1 1 0   1 1 0 1 1 1 1 1 1   1 1 1 0 1 1 1 0 1   1 1 1 0 1 1 1 0 0   1 1 1 0 1 1 0 1 1   1 1 1 0 1 1 0 1 0   1 1 1 0 1 1 0 0 1   1 1 1 0 1 1 0 0 0   1 1 1 0 1 0 1 1 1   1 1 1 0 1 0 1 1 0   1 1 1 0 1 0 1 0 1   1 1 1 0 1 0 1 0 0   1 1 1 0 1 0 0 1 1   1 1 1 0 1 0 0 1 0   1 1 1 0 1 0 0 0 1   1 1 1 0 1 0 0 0 0   1 1 1 0 0 1 1 1 1   1 1 1 0 0 1 1 1 0   1 1 1 0 0 1 1 0 1   1 1 1 0 0 1 1 0 0   1 1 1 0 0 1 0 1 1   1 1 1 0 0 1 0 1 0   1 1 1 0 0 1 0 0 1   1 1 1 0 0 1 0 0 0   1 1 1 0 0 0 1 1 1   1 1 1 0 0 0 1 1 0   1 1 1 0 0 0 1 0 1   1 1 1 0 0 0 1 0 0   1 1 1 0 0 0 0 1 1   1 1 1 0 0 0 0 1 0   1 1 1 0 0 0 0 0 1   1 1 1 0 0 0 0 0 0   1 1 0 1 1 1 1 1 0   1 1 0 1 1 1 1 0 1   1 1 0 1 1 1 1 0 0   1 1 0 1 1 1 0 1 1   1 1 0 1 1 1 0 0 1   1 1 0 1 1 1 0 0 0   1 1 0 1 1 0 1 1 1   1 1 0 1 1 0 1 1 0   1 1 0 1 1 0 1 0 1   1 1 0 1 1 0 1 0 0   1 1 0 1 1 0 0 1 1   1 1 0 1 1 0 0 1 0   1 1 0 1 1 0 0 0 1   1 1 0 1 1 0 0 0 0   1 1 0 1 0 1 1 1 1   1 1 0 1 0 1 1 1 0   1 1 0 1 0 1 1 0 1   1 1 0 1 0 1 1 0 0   1 1 0 1 0 1 0 1 1   1 1 0 1 0 1 0 1 0   1 1 0 1 0 1 0 0 1   1 1 0 1 0 1 0 0 1   1 1 0 1 0 1 0 0 0   1 1 0 1 0 0 1 1 1   1 1 0 1 0 0 1 1 0   1 1 0 1 0 0 1 0 1   1 1 0 1 0 0 1 0 0   1 1 0 1 0 0 0 1 1   1 1 0 1 0 0 0 1 0   1 1 0 1 0 0 0 0 0   1 1 0 1 0 0 0 0 0   1 1 0 0 1 1 1 1 1   1 1 0 0 1 1 1 1 0   1 1 0 0 1 1 1 0 1   1 1 0 0 1 1 1 0 0   1 1 0 0 1 1 0 1 1   1 1 0 0 1 1 0 1 0   1 1 0 0 1 1 0 0 1   1 1 0 0 1 1 0 0 0   1 1 0 0 1 0 1 1 1   1 1 0 0 1 0 1 1 0   1 1 0 0 1 0 1 0 1   1 1 0 0 1 0 1 0 0   1 1 0 0 1 0 0 1 1   1 1 0 0 1 0 0 1 0   1 1 0 0 1 0 0 0 1   1 1 0 0 1 0 0 0 0   1 1 0 0 0 1 1 1 1   1 1 0 0 0 1 1 1 0   1 1 0 0 0 1 1 0 1   1 1 0 0 0 1 1 0 0   1 1 0 0 0 1 0 1 1   1 1 0 0 0 1 0 1 0   1 1 0 0 0 1 0 0 1   1 1 0 0 0 0 1 0 0   1 1 0 0 0 0 0 1 1   1 1 0 0 0 0 0 1 0   1 1 0 0 0 0 0 0 1   1 1 0 0 0 0 0 0 0   1 0 1 1 1 1 1 1 0   1 0 1 1 1 1 1 0 1   1 0 1 1 1 1 1 0 0   1 0 1 1 1 1 0 1 1   1 0 1 1 1 1 0 1 0   1 0 1 1 1 1 0 0 1   1 0 1 1 1 1 0 0 0   1 0 1 1 1 0 1 1 1   1 0 1 1 1 0 1 1 0   1 0 1 1 1 0 1 0 1   1 0 1 1 1 0 1 0 0   1 0 1 1 1 0 0 1 1   1 0 1 1 1 0 0 1 0   1 0 1 1 1 0 0 0 1   1 0 1 1 1 0 0 0 0   1 0 1 1 0 1 1 1 1   1 0 1 1 0 1 1 1 0   1 0 1 1 0 1 1 0 1   1 0 1 1 0 1 1 0 0   1 0 1 1 0 1 0 1 1   1 0 1 1 0 1 0 1 0   1 0 1 1 0 1 0 0 1   1 0 1 1 0 1 0 0 0   1 0 1 1 0 0 1 1 1   1 0 1 1 0 0 1 1 0   1 0 1 1 0 0 1 0 1   1 0 1 1 0 0 1 0 0   1 0 1 1 0 0 0 1 1   1 0 1 1 0 0 0 1 0   1 0 1 1 0 0 0 0 1   1 0 1 1 0 0 0 0 0   1 0 1 0 1 1 1 1 1   1 0 1 0 1 1 1 0 1   1 0 1 0 1 1 1 0 0   1 0 1 0 1 1 0 1 1   1 0 1 0 1 1 0 1 0   1 0 1 0 1 1 0 0 1   1 0 1 0 1 1 0 0 0   1 0 1 0 1 0 1 1 1   1 0 1 0 1 0 1 1 0   1 0 1 0 1 0 1 0 1   1 0 1 0 1 0 1 0 1   1 0 1 0 1 0 0 1 1   1 0 1 0 1 0 0 1 0   1 0 1 0 1 0 0 0 1   1 0 1 0 1 0 0 0 0   1 0 1 0 0 1 1 1 1   1 0 1 0 0 1 1 1 0   1 0 1 0 0 1 1 0 1   1 0 1 0 0 1 1 0 0   1 0 1 0 0 1 0 1 1   1 0 1 0 0 1 0 1 0   1 0 1 0 0 1 0 0 1   1 0 1 0 0 1 0 0 0   1 0 1 0 0 0 1 1 1   1 0 1 0 0 0 1 1 0   1 0 1 0 0 0 1 0 1   1 0 1 0 0 0 1 0 0   1 0 1 0 0 0 0 1 1   1 0 1 0 0 0 0 1 0   1 0 1 0 0 0 0 0 1   1 0 1 0 0 0 0 0 0   1 0 0 1 1 1 1 1 0   1 0 0 1 1 1 1 0 1   1 0 0 1 1 1 1 0 0   1 0 0 1 1 1 0 1 1   1 0 0 1 1 1 0 1 0   1 0 1 1 1 0 0 1 0   1 0 1 1 1 0 0 0 1   1 0 1 1 1 0 0 0 0   1 0 1 1 0 1 1 1 1   1 0 1 1 0 1 1 1 0   1 0 1 1 0 1 1 0 1   1 0 1 1 0 1 1 0 0   1 0 1 1 0 1 0 1 1   1 0 1 1 0 1 0 1 0   1 0 1 1 0 1 0 0 1   1 0 1 1 0 1 0 0 0   1 0 1 1 0 0 1 1 1   1 0 1 1 0 0 1 1 0   1 0 1 1 0 1 0 0 1   1 0 1 1 0 1 0 0 0   1 0 1 1 0 0 1 1 1   1 0 1 1 0 0 1 1 0   1 0 1 1 0 0 1 0 1   1 0 1 1 0 0 1 0 0   1 0 1 1 0 0 0 1 1   1 0 1 1 0 0 0 1 0   1 0 1 1 0 0 0 0 1   1 0 1 1 0 0 0 0 0   1 0 1 0 1 1 1 1 1   1 0 1 0 1 1 1 0 1   1 0 1 0 1 1 1 0 0   1 0 1 0 1 1 0 1 1   1 0 1 0 1 1 0 1 0   1 0 1 0 1 1 0 0 1   1 0 1 0 1 1 0 0 0   1 0 1 0 1 0 1 1 1   1 0 1 0 1 0 1 1 0   1 0 1 0 1 0 1 0 1   1 0 1 0 1 0 1 0 0   1 0 1 0 1 0 0 1 1   1 0 1 0 1 0 0 1 0   1 0 1 0 1 0 0 0 1   1 0 1 0 1 0 0 0 0   1 0 1 0 0 1 1 1 1   1 0 1 0 0 1 1 1 0   1 0 1 0 0 1 1 0 1   1 0 1 0 0 1 1 0 0   1 0 1 0 0 1 0 1 1   1 0 1 0 0 1 0 1 0   1 0 1 0 0 1 0 0 1   1 0 1 0 0 1 0 0 0   1 0 1 0 0 0 1 1 1   1 0 1 0 0 0 1 1 0   1 0 1 0 0 0 1 0 1   1 0 1 0 0 0 1 0 0   1 0 1 0 0 0 0 1 1   1 0 1 0 0 0 0 1 0   1 0 1 0 0 0 0 0 1   1 0 1 0 0 0 0 0 0   1 0 0 1 1 1 1 1 1   1 0 0 1 1 1 1 1 0   1 0 0 1 1 1 1 0 1   1 0 0 1 1 1 1 1 0   1 0 0 1 1 1 1 0 1   1 0 0 1 1 1 1 0 0   1 0 0 1 1 1 0 1 1   1 0 0 1 1 1 0 1 0   1 0 0 1 1 1 0 0 1   1 0 0 1 1 1 0 0 0   1 0 0 1 1 0 1 1 1   1 0 0 1 1 0 1 1 0   1 0 0 1 1 0 1 0 1   1 0 0 1 1 0 1 0 0   1 0 0 1 1 0 0 1 1   1 0 0 1 1 0 0 1 0   1 0 0 1 1 0 0 0 1   1 0 0 1 1 0 0 0 0   1 0 0 1 0 1 1 1 1   1 0 0 1 0 1 1 1 0   1 0 0 1 0 1 1 0 1   1 0 0 1 0 1 1 0 0   1 0 0 1 0 1 0 1 1   1 0 0 1 0 1 0 1 0   1 0 0 1 0 1 0 0 1   1 0 0 1 0 1 0 0 0   1 0 0 1 0 0 1 1 1   1 0 0 1 0 0 1 1 0   1 0 0 1 0 0 1 0 1   1 0 0 1 0 0 1 0 0   1 0 0 1 0 0 0 1 1   1 0 0 1 0 0 0 1 0   1 0 0 1 0 0 0 0 1   1 0 0 1 0 0 0 0 0   1 0 0 0 1 1 1 1 1   1 0 0 0 1 1 1 1 0   1 0 0 0 1 1 1 0 1   1 0 0 0 1 1 1 0 0   1 0 0 0 1 1 0 1 1   1 0 0 0 1 1 0 1 0   1 0 0 0 1 1 0 0 1   1 0 0 0 1 1 0 0 0   1 0 0 0 1 0 1 1 1   1 0 0 0 1 0 1 1 0   1 0 0 0 1 0 1 0 1   1 0 0 0 1 0 1 0 0   1 0 0 0 1 0 0 1 1   1 0 0 0 1 0 0 1 0   1 0 0 0 1 0 0 0 1   1 0 0 0 1 0 0 0 0   1 0 0 0 0 1 1 1 1   1 0 0 0 0 0 1 1 0   1 0 0 0 0 0 1 0 1   1 0 0 0 0 0 1 0 0   1 0 0 0 0 0 0 1 1   1 0 0 0 0 0 0 1 0   1 0 0 0 0 0 0 0 1   1 0 0 0 0 0 0 0 0   0 1 1 1 1 1 1 1 0   0 1 1 1 1 1 1 0 1   0 1 1 1 1 1 1 0 0   0 1 1 1 1 1 0 1 1   0 1 1 1 1 1 0 1 0   0 1 1 1 1 1 0 0 1   0 1 1 1 1 1 0 0 0   0 1 1 1 1 0 1 1 1   0 1 1 1 1 0 1 1 0   0 1 1 1 1 0 1 0 1   0 1 1 1 1 0 1 0 0   0 1 1 1 1 0 0 1 1   0 1 1 1 1 0 0 1 0   0 1 1 1 1 0 0 0 1   0 1 1 1 1 0 0 0 0   0 1 1 1 0 1 1 1 1   0 1 1 1 0 1 1 0 0   0 1 1 1 0 1 0 1 1   0 1 1 1 0 1 0 1 0   0 1 1 1 0 1 0 0 1   0 1 1 1 0 1 0 0 0   0 1 1 1 0 0 1 1 1   0 1 1 1 0 0 1 1 0   0 1 1 1 0 0 1 0 1   0 1 1 1 0 0 1 0 0   0 1 1 1 0 0 0 1 1   0 1 1 1 0 0 0 1 0   0 1 1 1 0 0 0 0 1   0 1 1 1 0 0 0 0 0   0 1 1 0 1 1 1 1 0   0 1 1 0 1 1 1 0 1   0 1 1 0 1 1 1 0 0   0 1 1 0 1 1 0 1 1   0 1 1 0 1 1 0 1 0   0 1 1 0 1 1 0 0 1   0 1 1 0 1 1 0 0 0   0 1 1 0 1 0 1 1 1   0 1 1 0 1 0 1 1 0   0 1 1 0 1 0 1 0 1   0 1 1 0 1 0 0 1 0   0 1 1 0 1 0 0 0 1   0 1 1 0 1 0 0 0 0   0 1 1 0 0 1 1 1 1   0 1 1 0 0 1 1 1 0   0 1 1 0 0 1 1 0 1   0 1 1 0 0 1 1 0 0   0 1 1 0 0 1 0 1 1   0 1 1 0 0 1 0 1 0   0 1 1 0 0 1 0 0 1   0 1 1 0 0 1 0 0 0   0 1 1 0 0 0 1 1 1   0 1 1 0 0 0 1 1 0   0 1 1 0 0 0 1 0 1   0 1 1 0 0 0 1 0 0   0 1 1 0 0 0 0 1 1   0 1 1 0 0 0 0 1 0   0 1 1 0 0 0 0 0 1   0 1 1 0 0 0 0 0 0   0 1 0 1 1 1 1 1 0   0 1 0 1 1 1 1 0 1   0 1 0 1 1 1 1 0 0   0 1 0 1 1 1 0 1 1   0 1 0 1 1 1 0 1 0   0 1 0 1 1 1 0 0 1   0 1 0 1 1 1 0 0 0   0 1 0 1 1 0 1 1 1   0 1 0 1 1 0 1 1 0   0 1 0 1 1 0 1 0 1   0 1 0 1 1 0 1 0 0   0 1 0 1 1 0 0 1 1   0 1 0 1 1 0 0 1 0   0 1 0 1 1 0 0 0 1   0 1 0 1 1 0 0 0 0   0 1 0 1 0 1 1 1 1   0 1 0 1 0 1 1 1 0   0 1 0 1 0 1 1 0 1   0 1 0 1 0 1 1 0 0   0 1 0 1 0 1 0 1 1   0 1 0 1 0 1 0 1 0   0 1 0 1 0 1 0 0 1   0 1 0 1 0 1 0 0 0   0 1 0 1 0 1 0 0 0   0 1 0 1 0 0 1 1 1   0 1 0 1 0 0 1 1 0   0 1 0 1 0 0 1 0 1   0 1 0 1 0 0 1 0 0   0 1 0 1 0 0 0 1 1   0 1 0 1 0 0 0 1 0   0 1 0 1 0 0 0 0 1   0 1 0 1 0 0 0 0 0   0 1 0 0 1 1 1 1 1   0 1 0 0 1 1 1 1 0   0 1 0 0 1 1 1 0 1   0 1 0 0 1 1 1 0 0   0 1 0 0 1 1 0 1 1   0 1 0 0 1 1 0 1 0   0 1 0 0 1 1 0 0 1   0 1 0 0 1 1 0 0 0   0 1 0 0 1 0 1 1 1   0 1 0 0 1 0 1 1 0   0 1 0 0 1 0 1 0 1   0 1 0 0 1 0 1 0 0   0 1 0 0 1 0 0 1 1   0 1 0 0 1 0 0 1 0   0 1 0 0 1 0 0 0 1   0 1 0 0 1 0 0 0 0   0 1 0 0 0 1 1 1 1   0 1 0 0 0 1 1 1 0   0 1 0 0 0 1 1 0 1   0 1 0 0 0 1 1 0 0   0 1 0 0 0 1 0 1 1   0 1 0 0 0 1 0 1 0   0 1 0 0 0 1 0 0 1   0 1 0 0 0 1 0 0 0   0 1 0 0 0 0 1 1 1   0 1 0 0 0 0 1 1 0   0 1 0 0 0 0 1 0 1   0 1 0 0 0 0 1 0 0   0 1 0 0 0 0 0 1 1   0 1 0 0 0 0 0 0 1   0 1 0 0 0 0 0 0 0   0 0 1 1 1 1 1 1 1   0 0 1 1 1 1 1 1 0   0 0 1 1 1 1 1 0 1   0 0 1 1 1 1 1 0 0   0 0 1 1 1 1 0 1 1   0 0 1 1 1 1 0 1 0   0 0 1 1 1 1 0 0 1   0 0 1 1 1 1 0 0 0   0 0 1 1 1 0 1 1 1   0 0 1 1 1 0 1 1 0   0 0 1 1 1 0 1 0 1   0 0 1 1 1 0 1 0 0   0 0 1 1 1 0 0 1 1   0 0 1 1 1 0 0 0 1   0 0 1 1 1 0 0 0 0   0 0 1 1 0 1 1 1 1   0 0 1 1 0 1 1 1 0   0 0 1 1 0 1 1 0 1   0 0 1 1 0 1 1 0 0   0 0 1 1 0 1 0 1 1   0 0 1 1 0 1 0 1 0   0 0 1 1 0 1 0 0 1   0 0 1 1 0 1 0 0 0   0 0 1 1 0 0 1 1 1   0 0 1 1 0 0 1 1 0   0 0 1 1 0 0 1 0 1   0 0 1 1 0 0 1 0 0   0 0 1 1 0 0 0 1 1   0 0 1 1 0 0 0 1 0   0 0 1 1 0 0 0 0 1   0 0 1 0 1 1 1 1 1   0 0 1 0 1 1 1 1 0   0 0 1 0 1 1 1 0 1   0 0 1 0 1 1 1 0 0   0 0 1 0 1 0 1 1 0   0 0 1 0 1 0 1 0 1   0 0 1 0 1 0 1 0 0   0 0 1 0 1 0 0 1 1   0 0 1 0 1 0 0 1 0   0 0 1 0 1 0 0 0 1   0 0 1 0 1 0 0 0 0   0 0 1 0 0 1 1 1 1   0 0 1 0 0 1 1 1 0   0 0 1 0 0 1 1 0 1   0 0 1 0 0 1 1 0 0   0 1 0 0 0 1 0 1 1   0 0 1 0 0 1 0 0 0 1   0 0 0 1 1 1 1 1   0 0 0 1 1 1 1 1 1   0 0 0 0 1 1 1 1 1   0 0 0 0 1 1 1 1 0   0 0 0 0 1 1 1 0 1   0 0 0 0 1 1 1 0 0   0 0 0 0 1 1 0 1 1   0 0 0 0 1 1 0 1 0   0 0 0 0 1 1 0 0 1   0 0 0 0 1 1 0 0 0   0 0 0 0 1 0 1 1 1   0 0 0 0 1 0 1 1 0   0 0 0 0 1 0 0 0 1   0 0 0 0 1 0 0 0 0   0 0 0 0 0 1 1 1 1   0 0 0 0 0 1 1 1 0   0 0 0 0 0 1 1 0 1   0 0 0 0 0 1 1 0 0   0 0 0 0 0 1 0 1 1   0 0 0 0 0 1 0 1 0   0 0 0 0 0 1 0 0 1   0 0 0 0 0 1 0 0 0   0 0 0 0 0 0 1 1 1   0 0 0 0 0 0 1 1 0   0 0 0 0 0 0 1 0 1   0 0 0 0 0 0 1 0 0   0 0 0 0 0 0 0 1 1   0 0 0 0 0 0 0 1 0   0 0 0 0 0 0 0 0 1   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0 0   4 : 0 9   P M   2 0 2 4 - 1 2 - 2 6  
 1   2   1 0   1 1   1 2   2 0   2 1   2 2   1 0 0   1 0 1   1 0 2   1 1 0   1 1 1   1 1 2   1 2 0   1 2 1   1 2 2   2 0 0   2 0 1   2 0 2   2 1 0   2 1 1   2 1 2   2 2 1   2 2 2   1 0 0 0   1 0 0 2   1 0 1 0   1 0 1 1   1 0 2 1   1 0 2 2   1 1 0 0   1 1 0 1   1 1 0 2   1 1 1 0   1 1 1 1   1 1 1 2   1 1 2 0   1 1 2 1   1 1 2 2   1 2 0 1   1 2 0 2   1 2 1 0   1 2 1 1   1 2 1 2   1 2 2 1   1 2 2 2   2 0 0 0   2 0 0 1   2 0 0 2   2 0 1 0   2 0 1 1   2 0 1 2   2 0 2 0   2 0 2 1   2 0 2 2   2 1 0 0   2 1 0 1   2 1 0 2   2 1 1 0   2 1 1 1   2 1 1 2   2 1 2 0   2 1 2 1   2 1 2 2   2 2 0 0   2 2 0 1   2 2 0 2   2 2 1 0   2 2 1 1   2 2 1 2   2 2 2 0   2 2 2 1   2 2 2 2   1 0 0 0 0   1 0 0 0 1   1 0 0 0 2   1 0 0 1 0   1 0 0 1 1   1 0 0 1 2   1 0 0 2 0   1 0 0 2 1   1 0 0 2 2   1 0 1 0 0   1 0 1 0 1   1 0 1 0 2   1 0 1 1 0   1 0 1 1 1   1 0 1 1 2   1 0 1 2 0   1 0 1 2 1   1 0 1 2 2   1 0 2 0 0   1 0 2 0 1   1 0 2 0 2   1 0 2 1 0   1 0 2 1 1   1 0 2 1 2   1 0 2 2 0   1 0 2 2 1   1 0 2 2 2   1 1 0 0 0   1 1 0 0 1   1 1 0 0 2   1 1 0 1 0   1 1 0 1 1   1 1 0 1 2   1 1 0 2 0   1 1 0 2 1   1 1 0 2 2   1 1 1 0 0   1 1 1 0 1   1 1 1 0 2   1 1 1 1 0   1 1 1 1 1   1 1 1 1 2   1 1 1 2 0   1 1 1 2 1   1 1 1 2 2   1 1 2 0 0   1 1 2 0 1   1 1 2 0 2   1 1 2 1 0   1 1 2 1 1   1 1 2 1 2   1 1 2 2 0   1 1 2 2 1   1 1 2 2 2   1 2 0 0 0   1 2 0 0 1   1 2 0 0 2   1 2 0 1 0   1 2 0 1 1   1 2 0 1 2   1 2 0 2 0   1 2 0 2 1   1 2 0 2 2   1 2 1 0 0   1 2 1 0 1   1 2 1 0 2   1 2 1 1 0   1 2 1 1 1   1 2 1 1 2   1 2 1 2 0   1 2 1 2 1   1 2 1 2 2   1 2 2 0 0   1 2 2 0 1   1 2 2 0 2   1 2 2 1 0   1 2 2 1 1   1 2 2 1 2   1 2 2 2 0   1 2 2 2 1   1 2 2 2 2   2 0 0 0 0   2 0 0 0 1   2 0 0 0 2   2 0 0 1 0   2 0 0 1 1   2 0 0 1 2   2 0 0 2 0   2 0 0 2 1   2 0 0 2 2   2 0 1 0 0   2 0 1 0 1   2 0 1 0 2   2 0 1 1 0   2 0 1 1 1   2 0 1 1 2   2 0 1 2 0   2 0 1 2 1   2 0 1 2 2   2 0 2 0 0   2 0 2 0 1   2 0 2 0 2   2 0 2 1 0   2 0 2 1 1   2 0 2 1 2   2 0 2 2 0   2 0 2 2 1   2 0 2 2 2   2 1 0 0 0   2 1 0 0 1   2 1 0 0 2   2 1 0 1 0   2 1 0 1 1   2 1 0 1 2   2 1 0 2 0   2 1 0 2 1   2 1 0 2 2   2 1 1 0 0   2 1 1 0 1   2 1 1 0 2   2 1 1 1 0   2 1 1 1 1   2 1 1 1 2   2 1 1 2 0   2 1 1 2 1   2 1 1 2 2   2 1 2 0 0   2 1 2 0 1   2 1 2 0 2   2 1 2 1 0   2 1 2 1 1   2 1 2 1 2   2 1 2 2 0   2 1 2 2 1   2 1 2 2 2   2 2 0 0 0   2 2 0 0 1   2 2 0 0 2   2 2 0 1 0   2 2 0 1 1   2 2 0 1 2   2 2 0 2 0   2 2 0 2 1   2 2 0 2 2   2 2 1 0 0   2 2 1 0 1   2 2 1 0 2   2 2 1 1 0   2 2 1 1 1   2 2 1 1 2   2 2 1 2 0   2 2 1 2 1   2 2 1 2 2   2 2 2 0 0   2 2 2 0 1   2 2 2 0 2   2 2 2 1 0   2 2 2 1 1   2 2 2 1 2   2 2 2 2 0   2 2 2 2 1   2 2 2 2 2   1 0 0 0 0 0   1 0 0 0 0 1   1 0 0 0 0 2   1 0 0 0 1 0   1 0 0 0 1 1   1 0 0 0 1 2   1 0 0 0 2 0   1 0 0 0 2 1   1 0 0 0 2 2   1 0 0 1 0 0   1 0 0 1 0 1   1 0 0 1 0 2   1 0 0 1 1 0   1 0 0 1 1 1   1 0 0 1 1 2   1 0 0 1 2 0   1 0 0 1 2 1   1 0 0 1 2 2   1 0 0 2 0 0   1 0 0 2 0 1   1 0 0 2 0 2   1 0 0 2 1 0   1 0 0 2 1 1   1 0 0 2 1 2   1 0 0 2 2 0   1 0 0 2 2 1   1 0 0 2 2 2   1 0 1 0 0 0   1 0 1 0 0 1   1 0 1 0 0 2   1 0 1 0 1 0   1 0 1 0 1 1   1 0 1 0 1 2   1 0 1 0 2 0   1 0 1 0 2 1   1 0 1 0 2 2   1 0 1 1 0 0   1 0 1 1 0 1   1 0 1 1 0 2   1 0 1 1 1 0   1 0 1 1 1 1   1 0 1 1 1 2   1 0 1 1 2 0   1 0 1 1 2 1   1 0 1 1 2 2   1 0 1 2 0 0   1 0 1 2 0 1   1 0 1 2 0 2   1 0 1 2 1 0   1 0 1 2 1 0   1 0 1 2 1 1   1 0 1 2 1 2   1 0 1 2 2 0   1 0 1 2 2 1   1 0 1 2 2 2   1 0 2 0 0 0   1 0 2 0 0 1   1 0 2 0 0 2   1 0 2 0 1 0   1 0 2 0 1 1   1 0 2 0 1 2   1 0 2 0 2 0   1 0 2 0 2 1   1 0 2 0 2 2   1 0 2 1 0 0   1 0 2 1 0 1   1 0 2 1 0 2   1 0 2 1 1 0   1 0 2 1 1 1   1 0 2 1 2 0   1 0 2 1 2 1   1 0 2 1 2 2   1 0 2 2 0 0   1 0 2 2 0 1   1 0 2 2 0 2   1 0 2 2 1 0   1 0 2 2 1 1   1 0 2 2 1 2   1 0 2 2 2 0   1 0 2 2 2 1   1 0 2 2 2 2   1 1 0 0 0 0   1 1 0 0 0 1   1 1 0 0 0 2   1 1 0 0 1 0   1 1 0 0 1 1   1 1 0 0 1 2   1 1 0 0 2 0   1 1 0 0 2 1   1 1 0 0 2 2   1 1 0 1 0 0   1 1 0 1 0 1   1 1 0 1 0 2   1 1 0 1 1 0   1 1 0 1 1 1   1 1 0 1 1 2   1 1 0 1 2 0   1 1 0 1 2 1   1 1 0 1 2 2   1 1 0 2 0 0   1 1 0 2 0 1   1 1 0 2 0 2   1 1 0 2 1 0   1 1 0 2 1 1   1 1 0 2 1 2   1 1 0 2 2 0   1 1 0 2 2 1   1 1 0 2 2 2   1 1 1 0 0 0   1 1 1 0 0 0   1 1 1 0 0 1   1 1 1 0 0 2   1 1 1 0 1 0   1 1 1 0 1 1   1 1 1 0 1 2   1 1 1 0 2 0   1 1 1 0 2 1   1 1 1 0 2 2   1 1 1 1 0 0   1 1 1 1 0 2   1 1 1 1 1 0   1 1 1 1 1 1   1 1 1 1 1 2   1 1 1 1 2 0   1 1 1 1 2 1   1 1 1 1 2 2   1 1 1 2 0 0   1 1 1 2 0 1   1 1 1 2 0 2   1 1 1 2 1 0   1 1 1 2 1 1   1 1 1 2 1 2   1 1 1 2 2 0   1 1 1 2 2 1   1 1 1 2 2 2   1 1 2 0 0 0   1 1 2 0 0 1   1 1 2 0 0 2   1 1 2 0 1 0   1 1 2 0 1 1   1 1 2 0 1 2   1 1 2 0 2 0   1 1 2 0 2 1   1 1 2 0 2 2   1 1 2 1 0 0   1 1 2 1 0 1   1 1 2 1 0 2   1 1 2 1 1 0   1 1 2 1 1 1   1 1 2 1 2 0   1 1 2 1 2 1   1 1 2 1 2 2   1 1 2 2 0 0   1 1 2 2 0 1   1 1 2 2 0 2   1 1 2 2 1 0   1 1 2 2 1 1   1 1 2 2 1 2   1 1 2 2 2 0   1 1 2 2 2 1   1 1 2 2 2 2   1 2 0 0 0 0   1 2 0 0 0 1   1 2 0 0 0 2   1 2 0 0 1 0   1 2 0 0 1 1   1 2 0 0 1 2   1 2 0 0 2 0   1 2 0 0 2 1   1 2 0 0 2 2   1 2 0 1 0 0   1 2 0 1 0 1   1 2 0 1 0 2   1 2 0 1 1 0   1 2 0 1 1 1   1 2 0 1 1 2   1 2 0 1 2 0   1 2 0 1 2 1   1 2 0 1 2 2   1 2 0 2 0 0   1 2 0 2 0 1   1 2 0 2 0 2   1 2 0 2 1 0   1 2 0 2 1 1   1 2 0 2 1 2   1 2 0 2 2 0   1 2 0 2 2 1   1 2 0 2 2 2   1 2 1 0 0 0   1 2 1 0 0 1   1 2 1 0 0 2   1 2 1 0 1 0   1 2 1 0 1 1   1 2 1 0 1 2   1 2 1 0 2 0   1 2 1 0 2 1   1 2 1 0 2 2   1 2 1 1 0 0   1 2 1 1 0 1   1 2 1 1 0 2   1 2 1 1 1 0   1 2 1 1 1 1   1 2 1 1 1 2   1 2 1 1 2 0   1 2 1 1 2 1   1 2 1 1 2 2   1 2 1 2 0 0   1 2 1 2 0 1   1 2 1 2 0 2   1 2 1 2 1 0   1 2 1 2 1 1   1 2 1 2 1 2   1 2 1 2 2 0   1 2 1 2 2 1   1 2 1 2 2 2   1 2 2 0 0 0   1 2 2 0 0 1   1 2 2 0 0 2   1 2 2 0 1 0   1 2 2 0 1 1   1 2 2 0 1 2   1 2 2 0 2 0   1 2 2 0 2 1   1 2 2 0 2 2   1 2 2 1 0 0   1 2 2 1 0 1   1 2 2 1 0 2   1 2 2 1 1 0   1 2 2 1 1 1   1 2 2 1 1 2   1 2 2 1 2 0   1 2 2 1 2 1   1 2 2 1 2 2   1 2 2 2 2 0   1 2 2 2 0 0   1 2 2 2 0 1   1 2 2 2 0 2   1 2 2 2 1 0   1 2 2 2 1 1   1 2 2 2 1 2   1 2 2 2 2 0   1 2 2 2 2 1   1 2 2 2 2 2   2 0 0 0 0 0   2 0 0 0 0 1   2 0 0 0 0 2   2 0 0 0 1 0   2 0 0 0 1 1   2 0 0 0 1 2   2 0 0 0 2 0   2 0 0 0 2 1   2 0 0 0 2 2   2 0 0 1 0 0   2 0 0 1 0 1   2 0 0 1 0 2   2 0 0 1 1 0   2 0 0 1 1 1   2 0 0 1 2 0   2 0 0 1 2 1   2 0 0 1 2 2   2 0 0 2 0 0   2 0 0 2 0 1   2 0 0 2 0 2   2 0 0 2 1 0   2 0 0 2 1 1   2 0 0 2 1 2   2 0 0 2 2 0   2 0 0 2 2 1   2 0 0 2 2 2   2 0 1 0 0 0   2 0 1 0 0 1   2 0 1 0 0 2   2 0 1 0 1 0   2 0 1 0 1 1   2 0 1 0 1 2   2 0 1 0 2 0   2 0 1 0 2 1   2 0 1 0 2 2   2 0 1 1 0 0   2 0 1 1 0 1   2 0 1 1 0 2   2 0 1 1 1 0   2 0 1 1 1 1   2 0 1 1 1 2   2 0 1 1 2 0   2 0 1 1 2 1   2 0 1 1 2 2   2 0 1 2 0 0   2 0 1 2 1 0   2 0 1 2 0 1   2 0 1 2 0 2   2 0 1 2 1 0   2 0 1 2 1 1   2 0 1 2 1 2   2 0 1 2 2 0   2 0 1 2 2 1   2 0 1 2 2 2   2 0 2 0 0 0   2 0 2 0 0 1   2 0 2 0 0 2   2 0 2 0 1 0   2 0 2 0 1 1   2 0 2 0 1 2   2 0 2 0 2 0   2 0 2 0 2 1   2 0 2 0 2 2   2 0 2 1 0 0   2 0 2 1 0 1   2 0 2 1 0 2   2 0 2 1 1 0   2 0 2 1 1 1   2 0 2 1 1 2   2 0 2 1 2 0   2 0 2 1 2 1   2 0 2 1 2 2   2 0 2 2 0 0   2 0 2 2 0 1   2 0 2 2 0 2   2 0 2 2 1 0   2 0 2 2 1 1   2 0 2 2 1 2   2 0 2 2 2 0   2 0 2 2 2 1   2 0 2 2 2 2   2 1 0 0 0 0   2 1 0 0 0 1   2 1 0 0 0 2   2 1 0 0 1 0   2 1 0 0 1 1   2 1 0 0 1 2   2 1 0 0 2 0   2 1 0 0 2 1   2 1 0 0 2 2   2 1 0 1 0 0   2 1 0 1 0 1   2 1 0 1 0 2   2 1 0 1 1 0   2 1 0 1 1 1   2 1 0 1 1 2   2 1 0 1 2 0   2 1 0 1 2 1   2 1 0 1 2 2   2 1 0 2 0 0   2 1 0 2 0 1   2 1 0 2 0 2   2 1 0 2 1 0   2 1 0 2 1 1   2 1 0 2 1 2   2 1 0 2 2 0   2 1 0 2 2 1   2 1 0 2 2 2   2 1 1 0 0 0   2 1 1 0 0 1   2 1 1 0 0 2   2 1 1 0 1 0   2 1 1 0 1 1   2 1 1 0 1 2   2 1 1 0 2 0   2 1 1 0 2 1   2 1 1 0 2 2   2 1 1 1 0 0   2 1 1 1 0 1   2 1 1 1 0 2   2 1 1 1 1 0   2 1 1 1 1 1   2 1 1 1 2 0   2 1 1 1 2 1   2 1 1 1 2 2   2 1 1 2 0 0   2 1 1 2 0 1   2 1 1 2 0 2   2 1 1 2 1 0   2 1 1 2 1 1   2 1 1 2 1 2   2 1 1 2 2 0   2 1 1 2 2 1   2 1 1 2 2 2   2 1 2 0 0 0   2 1 2 0 0 1   2 1 2 0 0 2   2 1 2 0 1 0   2 1 2 0 1 1   2 1 2 0 1 2   2 1 2 0 2 0   2 1 2 0 2 1   2 1 2 0 2 2   2 1 2 1 0 0   2 1 2 1 0 1   2 1 2 1 0 2   2 1 2 1 1 0   2 1 2 1 1 1   2 1 2 1 1 2   2 1 2 1 2 0   2 1 2 1 2 1   2 1 2 1 2 2   2 1 2 2 0 0   2 1 2 2 0 1   2 1 2 2 0 2   2 1 2 2 1 0   2 1 2 2 1 1   2 1 2 2 1 2   2 1 2 2 1 2   2 1 2 2 2 0   2 1 2 2 2 1   2 1 2 2 2 2   2 2 0 0 0 0   2 2 0 0 0 1   2 2 0 0 0 2   2 2 0 0 1 0   2 2 0 0 1 1   2 2 0 0 1 2   2 2 0 0 2 0   2 2 0 0 2 1   2 2 0 0 2 2   2 2 0 1 0 0   2 2 0 1 0 1   2 2 0 1 0 2   2 2 0 1 1 0   2 2 0 1 1 1   2 2 0 1 1 2   2 2 0 1 2 0   2 2 0 1 2 1   2 2 0 1 2 2   2 2 0 2 0 0   2 2 0 2 0 1   2 2 0 2 0 2   2 2 0 2 1 0   2 2 0 2 1 2   2 2 0 2 1 1   2 2 0 2 1 2   2 2 0 2 2 0   2 2 0 2 2 1   2 2 0 2 2 2   2 2 1 0 0 0   2 2 1 0 0 1   2 2 1 0 0 2   2 2 1 0 1 0   2 2 1 0 1 1   2 2 1 0 1 2   2 2 1 0 2 0   2 2 1 0 2 1   2 2 1 1 0 0   2 2 1 1 0 0   2 2 1 1 0 1   2 2 1 1 0 2   2 2 1 1 1 0   2 2 1 1 1 1   2 2 1 1 1 2   2 2 1 1 2 0   2 2 1 1 2 1   2 2 1 1 2 2   2 2 1 2 0 0   2 2 1 2 0 1   2 2 1 2 0 2   2 2 1 2 1 0   2 2 1 2 1 1   2 2 1 2 1 2   2 2 1 2 2 0   2 2 1 2 2 1   2 2 1 2 2 2   2 2 0 0 0 0   2 2 2 0 0 0   2 2 2 0 0 1   2 2 2 0 0 2   2 2 2 0 1 0   2 2 2 0 1 1   2 2 2 0 1 2   2 2 2 0 2 0   2 2 2 0 2 1   2 2 2 0 2 2   2 2 2 1 0 0   2 2 2 1 0 1   2 2 2 1 0 2   2 2 2 1 1 0   2 2 2 1 1 1   2 2 2 1 1 2   2 2 2 1 2 0   2 2 2 1 2 1   2 2 2 1 2 2   2 2 2 2 0 0   2 2 2 2 0 1   2 2 2 2 0 2   2 2 2 2 1 0   2 2 2 2 1 1   2 2 2 2 1 2   2 2 2 2 2 0   2 2 2 2 2 1   2 2 2 2 2 2   1 0 0 0 0 0 0   1 0 0 0 0 0 1   1 0 0 0 0 2   1 0 0 0 0 1 0   1 0 0 0 0 1 1   1 0 0 0 0 1 2   1 0 0 0 0 2 0   1 0 0 0 0 2 1   1 0 0 0 0 2 2   1 0 0 0 1 0 0   1 0 0 0 1 0 1   1 0 0 0 1 0 2   1 0 0 0 1 1 0   1 0 0 0 1 1 1   1 0 0 0 1 1 2   1 0 0 0 1 2 0   1 0 0 0 1 2 1   1 0 0 0 1 2 2   1 0 0 0 2 0 0   1 0 0 0 2 0 1   1 0 0 0 2 0 2   1 0 0 0 2 1 0   1 0 0 0 2 1 1   1 0 0 0 2 1 2   1 0 0 0 2 2 0   1 0 0 0 2 2 1   1 0 0 0 2 2 2   1 0 0 1 0 0 0   1 0 0 1 0 0 1   1 0 0 1 0 0 2   1 0 0 1 0 1 0   1 0 0 1 0 1 1   1 0 0 1 0 1 2   1 0 0 1 0 2 0   1 0 0 1 0 2 1   1 0 0 1 0 2 2   1 0 0 1 1 0 0   1 0 0 1 1 0 1   1 0 0 1 1 0 2   1 0 0 1 1 1 0   1 0 0 1 1 1 1   1 0 0 1 1 1 2   1 0 0 1 1 2 0   1 0 0 1 1 2 1   1 0 0 1 1 2 2   1 0 0 1 2 0 0   1 0 0 1 2 0 1   1 0 0 1 2 0 2   1 0 0 1 2 1 0   1 0 0 1 2 1 1   1 0 0 1 2 1 2   1 0 0 1 2 2 0   1 0 0 1 2 2 1   1 0 0 1 2 2 2   1 0 0 2 0 0 0   1 0 0 2 0 0 1   1 0 0 2 0 0 2   1 0 0 2 0 1 0   1 0 0 2 0 1 1   1 0 0 2 0 1 2   1 0 0 2 0 2 0   1 0 0 2 0 2 1   1 0 0 2 0 2 2   1 0 0 2 1 0 0   1 0 0 2 1 0 1   1 0 0 2 1 0 2   1 0 0 2 1 1 0   1 0 0 2 1 1 1   1 0 0 2 1 1 2   1 0 0 2 1 2 0   1 0 0 2 1 2 1   1 0 0 2 1 2 2   1 0 0 2 2 0 0    
  
 4 : 2 3   P M   2 0 2 4 - 1 2 - 2 6  
  
 1 0 0 0 1 0 0 0   1 0 0 0 1 0 0 1   1 0 0 0 1 0 1 0   1 0 0 0 1 0 1 1   1 0 0 0 1 1 0 0   1 0 0 0 1 1 0 1   1 0 0 0 1 1 1 0   1 0 0 0 1 1 1 1   1 0 0 1 0 0 0 0   1 0 0 1 0 0 0 1   1 0 0 1 0 0 1 0   1 0 0 1 0 0 1 1   1 0 0 1 0 1 0 0   1 0 0 1 0 1 0 1   1 0 0 1 0 1 1 0   1 0 0 1 0 1 1 1   1 0 0 1 1 0 0 0   1 0 0 1 1 0 0 1   1 0 0 1 1 0 1 0   1 0 0 1 1 0 1 1   1 0 0 1 1 1 0 0   1 0 0 1 1 1 0 1   1 0 0 1 1 1 1 0   1 0 0 1 1 1 1 1   1 0 1 0 0 0 0 0   1 0 1 0 0 0 0 1   1 0 1 0 0 0 1 0   1 0 1 0 0 0 1 1   1 0 1 0 0 1 0 0   1 0 1 0 0 1 0 1   1 0 1 0 0 1 1 0   1 0 1 0 0 1 1 1   1 0 1 0 1 0 0 0   1 0 1 0 1 0 0 1   1 0 1 0 1 0 1 0   1 0 1 0 1 0 1 1   1 0 1 0 1 0 1 0   1 0 1 0 1 1 0 1   1 0 1 0 1 1 1 0   1 0 1 0 1 1 1 1   1 0 1 1 0 0 0 0   1 0 1 1 0 0 0 1   1 0 1 1 0 0 1 0   1 0 1 1 0 0 1 1   1 0 1 1 0 1 0 0   1 0 1 1 0 1 0 1   1 0 1 1 0 1 1 0   1 0 1 1 0 1 1 1   1 0 1 1 1 0 0 0   1 0 1 1 1 0 0 1   1 0 1 1 1 0 1 0   1 0 1 1 1 0 1 1   1 0 1 1 1 1 0 0   1 0 1 1 1 1 0 1   1 0 1 1 1 1 1 0   1 0 1 1 1 1 1 1   1 1 0 0 0 0 0 0   1 1 0 0 0 0 0 1   1 1 0 0 0 0 1 0   1 1 0 0 0 0 1 1   1 1 0 0 0 1 0 0   1 1 0 0 0 1 0 1   1 1 0 0 0 1 1 0   1 1 0 0 0 1 1 1   1 1 0 0 1 0 0 0   1 1 0 0 1 0 0 1   1 1 0 0 1 0 1 0   1 1 0 0 1 0 1 1   1 1 0 0 1 1 0 0   1 1 0 0 1 1 0 1   1 1 0 0 1 1 1 0   1 1 0 0 1 1 1 1   1 1 0 1 0 0 0 0   1 1 0 1 0 0 0 1   1 1 0 1 0 0 1 0   1 1 0 1 0 0 1 1   1 1 0 1 0 1 0 0   1 1 0 1 0 1 0 1   1 1 0 1 0 1 1 0   1 1 0 1 0 1 1 1   1 1 0 1 1 0 0 0   1 1 0 1 1 0 0 1   1 1 0 1 1 0 1 0   1 1 0 1 1 0 1 1   1 1 0 1 1 1 0 0   1 1 0 1 1 1 0 1   1 1 0 1 1 1 1 0   1 1 0 1 1 1 1 1   1 1 1 0 0 0 0 0   1 1 1 0 0 0 0 1   1 1 1 0 0 0 1 0   1 1 1 0 0 0 1 1   1 1 1 0 0 1 0 0   1 1 1 0 0 1 0 1   1 1 1 0 0 1 1 0   1 1 1 0 0 1 1 1   1 1 1 0 1 0 0 0   1 1 1 0 1 0 0 1   1 1 1 0 1 0 1 0   1 1 1 0 1 0 1 1   1 1 1 0 1 1 0 0   1 1 1 0 1 1 0 1   1 1 1 0 1 1 1 0   1 1 1 0 1 1 1 1   1 1 1 1 0 0 0 0   1 1 1 1 0 0 0 1   1 1 1 1 0 0 1 0   1 1 1 1 0 0 1 1   1 1 1 1 0 1 0 0   1 1 1 1 0 1 0 1   1 1 1 1 0 1 1 0   1 1 1 1 0 1 1 1   1 1 1 1 1 0 0 0   1 1 1 1 1 0 0 1   1 1 1 1 1 0 1 0   1 1 1 1 1 0 1 1   1 1 1 1 1 1 0 0   1 1 1 1 1 1 1 0   1 1 1 1 1 1 1 1   1 0 0 0 0 0 0 0 0   1 1 1 1 1 1 1 0   1 1 1 1 1 1 0 1   1 1 1 1 1 1 0 0   1 1 1 1 1 1 0 1   1 1 1 1 1 0 0 1   1 1 1 1 1 0 0 0   1 1 1 1 0 1 1 1   1 1 1 1 0 1 1 0   1 1 1 1 0 1 0 1   1 1 1 1 0 1 0 0   1 1 1 1 0 0 1 1   1 1 1 1 0 0 1 0   1 1 1 1 0 0 0 1   1 1 1 1 0 0 0 0   1 1 1 0 1 1 1 1   1 1 1 0 1 1 1 0   1 1 1 0 1 1 0 1   1 1 1 0 1 1 0 0   1 1 1 0 1 0 1 1   1 1 1 0 1 0 1 0   1 1 1 0 1 0 0 1   1 1 1 0 1 0 0 0   1 1 1 0 0 1 1 1   1 1 1 0 0 1 1 0   1 1 1 0 0 1 0 1   1 1 1 0 0 1 0 0   1 1 1 0 0 0 1 1   1 1 1 0 0 0 1 0   1 1 1 0 0 0 0 1   1 1 1 0 0 0 0 0   1 1 0 1 1 1 1 1   1 1 0 1 1 1 1 0   1 1 0 1 1 1 0 1   1 1 0 1 1 1 0 0   1 1 0 1 1 0 1 1   1 1 0 1 1 0 1 0   1 1 0 1 1 0 0 1   1 1 0 1 1 0 0 0   1 1 0 1 0 1 1 1   1 1 0 1 0 1 1 0   1 1 0 1 0 1 0 1   1 1 0 1 0 1 0 0   1 1 0 1 0 0 1 1   1 1 0 1 0 0 1 0   1 1 0 1 0 0 0 1   1 1 0 1 0 0 0 0   1 1 0 0 1 1 1 1   1 1 0 0 1 1 1 0   1 1 0 0 1 1 0 1   1 1 0 0 1 1 0 0   1 1 0 0 1 0 1 1   1 1 0 0 1 0 1 0   1 1 0 0 1 0 0 1   1 1 0 0 1 0 0 0   1 1 0 0 0 1 1 1   1 1 0 0 0 1 1 0   1 1 0 0 0 1 0 1   1 1 0 0 0 1 0 0   1 1 0 0 0 0 1 1   1 1 0 0 0 0 1 0   1 1 0 0 0 0 0 1   1 1 0 0 0 0 0 0   1 0 1 1 1 1 1 0   1 0 1 1 1 0 1 1   1 0 1 1 1 0 1 0   1 0 1 1 1 0 0 1   1 0 1 1 1 0 0 0   1 0 1 1 0 1 1 1   1 0 1 1 0 1 1 0   1 0 1 1 0 1 0 1   1 0 1 1 0 1 0 0   1 0 1 1 0 0 1 1   1 0 1 1 0 0 0 1   1 0 1 1 0 0 0 0   1 0 1 0 1 1 1 1   1 0 1 0 1 1 1 0   1 0 1 0 1 1 0 1   1 0 1 0 1 1 0 0   1 0 1 0 1 0 1 1   1 0 1 0 1 0 1 0   1 0 1 0 1 0 0 1   1 0 1 0 1 0 0 0   1 0 1 0 1 0 0 1   1 0 1 0 1 0 0 0   1 0 1 0 0 1 1 1   1 0 1 0 0 1 1 0   1 0 1 0 0 1 0 1   1 0 1 0 0 1 0 0   1 0 1 0 0 0 1 1   1 0 1 0 0 0 1 0   1 0 1 0 0 0 0 1   1 0 1 0 0 0 0 0   1 0 0 1 1 1 1 1   1 0 0 0 1 1 1 0   1 0 0 0 1 1 1 0   1 0 0 0 1 1 0 0   1 0 0 0 1 0 1 1   1 0 0 0 1 0 1 1   1 0 0 0 1 0 1 0   1 0 0 0 1 0 0 1   1 0 0 0 1 0 0 0   1 0 0 0 0 0 1 1   1 0 0 0 0 0 1 1   1 0 0 0 0 0 1 0   1 0 0 0 0 0 0 1   1 0 0 0 0 0 0 0   0 1 1 1 1 1 1 0   0 1 1 1 1 1 0 1   0 1 1 1 1 1 0 0   0 1 1 1 1 0 1 1   0 1 1 1 1 0 1 0   0 1 1 1 1 0 0 1   0 1 1 1 1 0 0 0   0 1 1 1 0 1 1 1   0 1 1 1 0 1 1 0   0 1 1 1 0 1 0 1   0 1 1 1 0 1 0 0   0 1 1 1 0 0 1 1   0 1 1 1 0 0 1 0   0 1 1 1 0 0 0 1   0 1 1 1 0 0 0 0   0 1 1 0 1 1 1 1   0 1 1 0 1 1 1 0   0 1 1 0 1 1 0 1   0 1 1 0 1 1 0 0   0 1 1 0 1 0 1 1   0 1 1 0 1 0 1 0   0 1 1 0 1 0 0 1   0 1 1 0 1 0 0 0   0 1 1 0 0 1 1 1   0 1 1 0 0 1 1 0   0 1 1 0 0 1 0 1   0 1 1 0 0 1 0 0   0 1 1 0 0 0 1 1   0 1 1 0 0 0 1 0   0 1 1 0 0 0 0 1   0 1 1 0 0 0 0 0   0 1 0 1 1 1 1 0   0 1 0 1 1 1 0 1   0 1 0 1 1 1 0 0   0 1 0 1 1 0 1 1   0 1 0 1 1 0 1 0   0 1 0 1 1 0 0 1   0 1 0 1 1 0 0 0   0 1 0 1 0 1 1 1   0 1 0 1 0 1 1 0   0 1 0 1 0 1 0 1   0 1 0 1 0 1 0 0   0 1 0 1 0 0 1 1   0 1 0 1 0 0 1 0   0 1 0 1 0 0 0 1   0 1 0 1 0 0 0 0   0 1 0 0 1 1 1 1   0 1 0 0 1 1 1 0   0 1 0 0 1 1 0 1   0 1 0 0 1 1 0 0   0 1 0 0 1 0 1 1   0 1 0 0 1 0 1 0   0 1 0 0 1 0 0 1   0 1 0 0 1 0 0 0   0 1 0 0 0 1 1 1   0 1 0 0 0 1 1 0   0 1 0 0 0 1 0 1   0 1 0 0 0 1 0 0   0 1 0 0 0 0 1 1   0 1 0 0 0 0 1 0   0 1 0 0 0 0 0 1   0 1 0 0 0 0 0 0   0 0 1 1 1 1 1 1   0 0 1 1 1 1 1 0   0 0 1 1 1 1 0 1   0 0 1 1 1 1 0 0   0 0 1 1 1 0 1 1   0 0 1 1 1 0 1 0   0 0 1 1 1 0 0 1   0 0 1 1 1 0 0 0   0 0 1 1 0 1 1 1   0 0 1 1 0 1 1 0   0 0 1 1 0 1 0 1   0 0 1 1 0 0 1 1   0 0 1 1 0 0 1 0   0 0 1 1 0 0 0 1   0 0 1 1 0 0 0 0   0 0 1 0 1 1 1 1   0 0 1 0 1 1 1 0   0 0 1 0 1 1 0 1   0 0 1 0 1 1 0 0   0 0 1 0 1 0 1 1   0 0 1 0 1 0 1 0   0 0 1 0 1 0 0 1   0 0 1 0 1 0 0 0   0 0 1 0 0 1 1 1   0 0 1 0 0 1 1 0   0 0 1 0 0 1 0 1   0 0 1 0 0 1 0 0   0 0 1 0 0 0 1 1   0 0 1 0 0 0 1 0   0 0 1 0 0 0 0 1   0 0 1 0 0 0 0 0   0 0 0 1 1 1 1 0   0 0 0 1 1 1 0 1   0 0 0 1 1 1 0 0   0 0 0 1 1 0 1 1   0 0 0 1 1 0 1 0   0 0 0 1 1 0 0 1   0 0 0 1 1 0 0 0   0 0 0 1 0 1 1 1   0 0 0 1 0 1 1 0   0 0 0 1 0 1 1 0   0 0 0 1 0 1 0 1   0 0 0 1 0 1 0 0   0 0 0 1 0 0 1 1   0 0 0 1 0 0 1 0   0 0 0 1 0 0 0 1   0 0 0 1 0 0 0 0   0 0 0 0 1 1 1 1   0 0 0 0 1 1 1 0   0 0 0 0 1 1 0 1   0 0 0 0 1 1 0 0   0 0 0 0 1 0 1 1   0 0 0 0 1 0 1 0   0 0 0 0 1 0 0 1   0 0 0 0 1 0 0 0   0 0 0 0 0 1 1 1   0 0 0 0 0 1 1 0   0 0 0 0 0 1 1 0   0 0 0 0 0 1 0 1   0 0 0 0 0 1 0 0   0 0 0 0 0 0 1 1   0 0 0 0 0 0 0 1   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   0 0 0 0 0 0 0 0   4 : 3 3   P M   2 0 2 4 - 1 2 - 2 6  
  
 1 0 0   4   1 0 1   1 1 0   1 1 1   1 0 0 0   1 0 0 1   1 0 1 0   1 0 1 1   1 1 0 0   1 1 0 1   1 1 1 0   1 1 1 1   1 0 0 0 0   1 0 0 0 1   1 0 0 1 0   1 0 0 1 1   1 0 1 0 0   1 0 1 0 1   1 0 1 1 0   1 0 1 1 1   1 1 0 0 0   1 1 0 0 1   1 1 0 1 0   1 1 0 1 1   1 1 1 0 0   1 1 1 0 1   1 1 1 1 0   1 1 1 1 1   1 0 0 0 0 0   1 0 0 0 0 1   1 0 0 0 1 0   1 0 0 0 1 1   1 0 0 1 0 0   1 0 0 1 0 1   1 0 0 1 1 0   1 0 0 1 1 1   1 0 1 0 0 0   1 0 1 0 0 1   1 0 1 0 1 0   1 0 1 0 1 1   1 0 1 1 0 0   1 0 1 1 0 1   1 0 1 1 1 0   1 0 1 1 1 1   1 1 0 0 0 0   1 1 0 0 0 1   1 1 0 0 1 0   1 1 0 0 1 1   1 1 0 1 0 0   1 1 0 1 0 1   1 1 0 1 1 0   1 1 0 1 1 1   1 1 1 0 0 0   1 1 1 0 0 1   1 1 1 0 0 1   1 1 1 0 1 0   1 1 1 0 1 1   1 1 1 1 0 0   1 1 1 1 0 1   1 1 1 1 1 0   1 1 1 1 1 1   1 0 0 0 0 0 0   1 1 1 1 1 1   1 1 1 1 1 0   1 1 1 1 0 1   1 1 1 1 0 0   1 1 1 0 1 1   1 1 1 0 1 0   1 1 1 0 0 1   1 1 1 0 0 0   1 1 0 1 1 1   1 1 0 1 1 0   1 1 0 1 0 1   1 1 0 1 0 0   1 1 0 0 1 1   1 1 0 0 1 0   1 1 0 0 0 1   1 1 0 0 0 0   1 0 1 1 1 1   1 0 1 1 1 0   1 0 1 1 0 1   1 0 1 1 0 0   1 0 1 0 1 1   1 0 1 0 1 0   1 0 1 0 0 1   1 0 1 0 0 0   1 0 0 1 1 1   1 0 0 1 1 0   1 0 0 1 0 1   1 0 0 1 0 0   1 0 0 0 1 1   1 0 0 0 1 0   1 0 0 0 0 1   1 0 0 0 0 0   1 1 1 1 1   1 1 1 1 0   1 1 1 0 1   1 1 1 0 0   1 1 0 1 1   1 1 0 1 0   1 1 0 0 1   1 1 0 0 0   1 0 1 1 1   1 0 1 1 0   1 0 1 0 1   1 0 1 0 0   1 0 0 1 1   1 0 0 1 0   1 0 0 0 1   1 0 0 0 0   1 1 1 1   1 1 1 0   1 1 0 1   1 1 0 0   1 0 1 1   1 0 1 0   1 0 0 1   1 0 0 0   1 1 1   1 1 0   1 0 1   1 0 0   1 1   1 0   1   0   + =   1   = =   1   + =   1 0   1 1   1 0 0   1 0 1   1 1 0   1 1 1   0 1 0 0   1 0 0 0   1 0 0 1   1 0 1 0   1 0 1 1   1 0 0 0 0   1 0 0 0 1   1 0 0 1 0   1 0 0 1 1   1 0 1 0 0   1 0 1 0 1   1 0 1 1 0   1 0 1 1 1   1 1 0 0 0   1 1 0 0 1   1 1 0 0 1   1 1 0 1 0   1 1 0 1 1   1 1 1 0 0   1 1 1 0 1   1 1 1 1 0   1 1 1 1 1   1 0 0 0 0 0   1 0 0 0 0 1   1 0 0 0 1 0   1 0 0 0 1 1   1 0 0 1 0 0   1 0 0 1 0 1   1 0 0 1 1 0   1 0 0 1 1 1   1 0 1 0 0 0   1 0 1 0 0 1   1 0 1 0 1 0   1 0 1 0 1 1   1 0 1 1 0 0   1 0 1 1 0 1   1 0 1 1 1 0   1 0 1 1 1 1   1 1 0 0 0 0   1 1 0 0 0 1   1 1 0 0 1 0   1 1 0 0 1 1   1 1 0 1 0 0   1 1 0 1 0 1   1 1 0 1 1 0   1 1 0 1 1 1   1 1 1 0 0 0   1 1 1 0 0 1   1 1 1 0 1 0   1 1 1 0 1 1   1 1 1 1 0 0   1 1 1 1 0 1   1 1 1 1 1 0   1 1 1 1 1 1   1 0 0 0 0 0 0   1 0 0 0 1 0 0 0   1 0 0 0 1 0 0 1   1 0 0 0 1 0 1 0   1 0 0 0 1 0 1 1   1 0 0 0 1 1 0 0   1 0 0 0 1 1 0 1   1 0 0 0 1 1 1 0   1 0 0 0 1 1 1   1 0 0 1 0 0 0   1 0 0 1 0 0 1   1 0 0 1 0 1 0   1 0 0 1 0 1 1   1 0 0 1 1 0 0   1 0 0 1 1 0 1   1 0 0 1 1 1 0   1 0 0 1 1 1 1   1 0 1 0 0 0 0   1 0 1 0 0 0 1   1 0 1 0 0 1 0   1 0 1 0 0 1 1   1 0 1 0 1 0 0   1 0 1 0 1 0 1   1 0 1 0 1 1 0   1 0 1 0 1 1 1   1 0 1 1 0 0 0   1 0 1 1 0 0 1   1 0 1 1 0 1 0   1 0 1 1 0 1 1   1 0 1 1 1 0 0   1 0 1 1 1 0 1   1 0 1 1 1 1 0   1 0 1 1 1 1 1   1 1 0 0 0 0   1 1 0 0 0 0 1   1 1 0 0 0 1 0   1 1 0 0 0 1 1   1 1 0 0 1 0 0   1 1 0 0 1 0 1   1 1 0 0 1 1 0   1 1 0 0 1 1 1   1 1 0 1 0 0 0   1 1 0 1 0 0 1   1 1 0 1 0 1 0   1 1 0 1 0 1 1   1 1 0 1 1 0 0   1 1 0 1 1 0 1   1 1 0 1 1 1 0   1 1 0 1 1 1 1   1 1 1 0 0 0 0   1 1 1 0 0 0 1   1 1 1 0 0 1 0   1 1 1 0 0 1 1   1 1 1 0 1 0 0   1 1 1 0 1 0 1   1 1 1 0 1 1 0   1 1 1 0 1 1 1   1 1 1 1 0 0 0   1 1 1 1 0 0 1   1 1 1 1 0 1 0   1 1 1 1 0 1 1   1 1 1 1 1 0 0   1 1 1 1 1 0 1   1 1 1 1 1 1 0   1 1 1 1 1 1 1   1 0 0 0 0 0 0 0   1 0 0 0 0 0 0 1   1 0 0 0 1 0 0 0   1 0 0 0 1 0 0 1   1 0 0 0 1 0 1 0   1 0 0 0 1 0 1 1   1 0 0 0 1 1 0 0   1 0 0 1 1 0 1   1 0 0 0 1 1 1 0   1 0 0 0 1 1 1 1   1 0 0 1 0 0 0 0   1 0 0 1 0 0 0 1   1 0 0 1 0 0 1 0   1 0 0 1 0 0 1 1   1 0 0 1 0 1 0 0   1 0 0 1 0 1 0 1   1 0 0 1 0 1 1 0   1 0 0 1 0 1 1 1   1 0 0 1 1 0 0 0   1 0 0 1 1 0 0 1   1 0 0 1 1 0 1 0   1 0 0 1 1 0 1 1   1 0 0 1 1 1 0 0   1 0 0 1 1 1 0 1   1 0 0 1 1 1 1 0   1 0 0 1 1 1 1 1   1 0 1 0 0 0 0 0   1 0 1 0 0 0 0 1   1 0 1 0 0 0 1 0   1 0 1 0 0 0 1 1   1 0 1 0 0 1 0 0   1 0 1 0 0 1 0 1   1 0 1 0 0 1 1 0   1 0 1 0 0 1 1 1   1 0 1 0 1 0 0 0   1 0 1 0 1 0 0 1   1 0 1 0 1 0 1 0   1 0 1 0 1 0 1 1   1 0 1 0 1 1 0 0   1 0 1 0 1 1 0 1   1 0 1 0 1 1 1 0   1 0 1 0 1 1 1 1   1 0 1 1 0 0 0 0   1 0 1 1 0 0 0 1   1 0 1 1 0 0 1 0   1 0 1 1 0 0 1 1   1 0 1 1 0 1 0 0   1 0 1 1 0 1 0 1   1 0 1 1 0 1 1 0   1 0 1 1 0 1 1 1   1 0 1 1 1 0 0 0   1 0 1 1 1 0 0 1   1 0 1 1 1 0 0 1   1 0 1 1 1 0 0 1   1 0 1 1 1 0 1 0   1 0 1 1 1 0 1 1   1 0 1 1 1 1 0 0   1 0 1 1 1 1 0 1   1 0 1 1 1 1 1 0   1 0 1 1 1 1 1   1 1 0 0 0 0 0 0   1 1 0 0 0 0 0 1   1 1 0 0 0 0 1 0   1 1 0 0 0 0 1 1   1 1 0 0 0 1 0 0   1 1 0 0 0 1 0 1   1 1 0 0 0 1 1 0   1 1 0 0 0 1 1 1   1 1 0 0 1 0 0 0   1 1 0 0 1 0 0 1   1 1 0 0 1 0 1 0   1 1 0 0 1 0 1 1   1 1 0 0 1 1 0 0   1 1 0 0 1 1 1 0   1 1 0 0 1 1 1 1   1 1 0 1 0 0 0 0   1 1 0 1 0 0 0 1   1 1 0 1 0 0 1 0   1 1 0 1 0 0 1 1   1 1 0 1 0 1 0 0   1 1 0 1 0 1 0 1   1 1 0 1 0 1 1 0   1 1 0 1 0 1 1 1   1 1 0 1 1 0 0 0   1 1 0 1 1 0 0 1   1 1 0 1 1 0 1 0   1 1 0 1 1 0 1 1   1 1 0 1 1 1 0 0   1 1 0 1 1 1 0 1   1 1 0 1 1 1 1 0   1 1 0 1 1 1 1 1   1 1 1 0 0 0 0 0   1 1 1 0 0 0 0 1   1 1 1 0 0 0 1 0   1 1 1 0 0 0 1 1   1 1 1 0 0 1 0 0   1 1 1 0 0 1 0 1   1 1 1 0 0 1 1 0   1 1 1 0 0 1 1 1   1 1 1 0 1 0 0 0   1 1 1 0 1 0 0 1   1 1 1 0 1 0 1 0   1 1 1 0 1 0 1 1   1 1 1 0 1 1 0 0   1 1 1 0 1 1 0 1   1 1 1 0 1 1 1 0   1 1 1 0 1 1 1   1 1 1 1 0 0 0 0   1 1 1 1 0 0 0 1   1 1 1 1 0 0 1 0   1 1 1 1 0 0 1 1   1 1 1 1 0 1 0 0   1 1 1 1 0 1 0 1   1 1 1 1 0 1 1 0   1 1 1 1 0 1 1 1   1 1 1 1 1 0 0 0   1 1 1 1 1 0 1 0   1 1 1 1 1 0 1 0   1 1 1 1 1 0 1 1   1 1 1 1 1 1 0 0   1 1 1 1 1 1 0 1   1 1 1 1 1 1 1 0   1 1 1 1 1 1 1 1   1 1 1 1 1 1 1 0   1 1 1 1 1 1 0 1   1 1 1 1 1 1 0 0   1 1 1 1 1 0 1 1   1 1 1 1 1 0 1 0   1 1 1 1 1 0 0 1   1 1 1 1 1 0 0 0   1 1 1 1 0 0 0 0  
  
 4 : 4 4   P M   2 0 2 4 - 1 2 - 2 6  
 